/*
* Copyright 2018 ARDUINO SA (http://www.arduino.cc/)
* This file is part of Vidor IP.
* Copyright (c) 2018
* Authors: Dario Pennisi
*
* This software is released under:
* The GNU General Public License, which covers the main part of 
* Vidor IP
* The terms of this license can be found at:
* https://www.gnu.org/licenses/gpl-3.0.en.html
*
* You can be released from the requirements of the above licenses by purchasing
* a commercial license. Buying such a license is mandatory if you want to modify or
* otherwise use the software for commercial activities involving the Arduino
* software without disclosing the source code of your own applications. To purchase
* a commercial license, send an email to license@arduino.cc.
*
*/

module MKRVIDOR4000_top
(
  // system signals
  input         iCLK,
  input         iRESETn,
  input         iSAM_INT,
  output        oSAM_INT,
  
  // SDRAM
  output        oSDRAM_CLK,
  output [11:0] oSDRAM_ADDR,
  output [1:0]  oSDRAM_BA,
  output        oSDRAM_CASn,
  output        oSDRAM_CKE,
  output        oSDRAM_CSn,
  inout  [15:0] bSDRAM_DQ,
  output [1:0]  oSDRAM_DQM,
  output        oSDRAM_RASn,
  output        oSDRAM_WEn,

  // SAM D21 PINS
  inout         bMKR_AREF,
  inout  [6:0]  bMKR_A,
  inout  [14:0] bMKR_D,
  
  // Mini PCIe
  inout         bPEX_RST,
  inout         bPEX_PIN6,
  inout         bPEX_PIN8,
  inout         bPEX_PIN10,
  input         iPEX_PIN11,
  inout         bPEX_PIN12,
  input         iPEX_PIN13,
  inout         bPEX_PIN14,
  inout         bPEX_PIN16,
  inout         bPEX_PIN20,
  input         iPEX_PIN23,
  input         iPEX_PIN25,
  inout         bPEX_PIN28,
  inout         bPEX_PIN30,
  input         iPEX_PIN31,
  inout         bPEX_PIN32,
  input         iPEX_PIN33,
  inout         bPEX_PIN42,
  inout         bPEX_PIN44,
  inout         bPEX_PIN45,
  inout         bPEX_PIN46,
  inout         bPEX_PIN47,
  inout         bPEX_PIN48,
  inout         bPEX_PIN49,
  inout         bPEX_PIN51,

  // NINA interface
  inout         bWM_PIO1,
  inout         bWM_PIO2,
  inout         bWM_PIO3,
  inout         bWM_PIO4,
  inout         bWM_PIO5,
  inout         bWM_PIO7,
  inout         bWM_PIO8,
  inout         bWM_PIO18,
  inout         bWM_PIO20,
  inout         bWM_PIO21,
  inout         bWM_PIO27,
  inout         bWM_PIO28,
  inout         bWM_PIO29,
  inout         bWM_PIO31,
  input         iWM_PIO32,
  inout         bWM_PIO34,
  inout         bWM_PIO35,
  inout         bWM_PIO36,
  input         iWM_TX,
  inout         oWM_RX,
  inout         oWM_RESET,

  // HDMI output
  output [2:0]  oHDMI_TX,
  output        oHDMI_CLK,

  inout         bHDMI_SDA,
  inout         bHDMI_SCL,
  
  input         iHDMI_HPD,
  
  // MIPI input
  input  [1:0]  iMIPI_D,
  input         iMIPI_CLK,
  inout         bMIPI_SDA,
  inout         bMIPI_SCL,
  inout  [1:0]  bMIPI_GP,

  // Q-SPI Flash interface
  output        oFLASH_SCK,
  output        oFLASH_CS,
  inout         oFLASH_MOSI,
  inout         iFLASH_MISO,
  inout         oFLASH_HOLD,
  inout         oFLASH_WP

);

// signal declaration

wire        wOSC_CLK;

wire        wCLK8,wCLK24, wCLK64, wCLK120;

wire [31:0] wJTAG_ADDRESS, wJTAG_READ_DATA, wJTAG_WRITE_DATA, wDPRAM_READ_DATA;
wire        wJTAG_READ, wJTAG_WRITE, wJTAG_WAIT_REQUEST, wJTAG_READ_DATAVALID;
wire [4:0]  wJTAG_BURST_COUNT;
wire        wDPRAM_CS;

wire [7:0]  wDVI_RED,wDVI_GRN,wDVI_BLU;
wire        wDVI_HS, wDVI_VS, wDVI_DE;

wire        wVID_CLK, wVID_CLKx5;
wire        wMEM_CLK;

assign wVID_CLK   = wCLK24;
assign wVID_CLKx5 = wCLK120;
assign wCLK8      = iCLK;

// internal oscillator
cyclone10lp_oscillator   osc
  ( 
  .clkout(wOSC_CLK),
  .oscena(1'b1));

// system PLL
SYSTEM_PLL PLL_inst(
  .areset(1'b0),
  .inclk0(wCLK8),
  .c0(wCLK24),
  .c1(wCLK120),
  .c2(wMEM_CLK),
  .c3(oSDRAM_CLK),
  .c4(wFLASH_CLK),
  .locked()
  );
  

wire [10:0]  aa, tt;  // GL-25jan2023
wire         by, as, ts, c1, c2, tr, sm1, sm2, st, go;

// D0 generated by CPU (User type G)

Schema Schema_inst
(
.F36MHz(wOSC_CLK),    // Main Clock

.MKR_D0(bMKR_D[0]),   // Tshift to CPU

.MKR_D1(bMKR_D[1]),   // INPUT  channel 1 with Trigger
.MKR_D2(bMKR_D[2]),   // INPUT  channel 2
.MKR_D3(bMKR_D[3]),
.MKR_D4(bMKR_D[4]),
.MKR_D5(bMKR_D[5]),
.MKR_D6(bMKR_D[6]),
.MKR_D7(bMKR_D[7]),   // INPUT  channel 7
.MKR_D8(bMKR_D[8]),   // OUTPUT channel 1
.MKR_D9(bMKR_D[9]),
.MKR_D10(bMKR_D[10]),
.MKR_D11(bMKR_D[11]),
.MKR_D12(bMKR_D[12]),
.MKR_D13(bMKR_D[13]),
.MKR_D14(bMKR_D[14]), // OUTPUT channel 7

//     (bMKR_A[0]) used by CPU to generate signal

.MKR_A1(bMKR_A[1]),   // ByAV to CPU 

.MKR_A2(bMKR_A[2]),   // Latch
.MKR_A3(bMKR_A[3]),   // Reset
.MKR_A4(bMKR_A[4]),   // Clk

.iByAv(by),
.iAshift(as),
.iTshift(ts),
.iClr1(c1),
.iClr2(c2),

.oSM1clk(sm1),
.oSM2clk(sm2),
.oTrigger(tr),
.A(aa),
.T(tt)
);

SM1 SM1_inst
(
.reset(),
.iSM1clk(sm1),
.iTrigger(tr),
.A(aa),
.iA5(bMKR_A[5]),    //    generated by CPU
.iA6(bMKR_A[6]),    //    generated by CPU
.iGO(go),

.oAshift(as),		  // Acquisition shift
.oClr1(c1),			  // Clear counters
.oStart(st)         // Start SM2
);

SM2 SM2_inst
(
.reset(),
.iSM2clk(sm2),
.T(tt),
.iStart(st),

.oByAv(by),
.oTshift(ts),		  // Transfer shift
.oClr2(c2),			  // Clear counters
.oGo(go)
);

reg [5:0] rRESETCNT;

always @(posedge wMEM_CLK)
begin
  if (!rRESETCNT[5])
  begin
  rRESETCNT<=rRESETCNT+1;
  end
end

endmodule
